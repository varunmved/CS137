//adder.v 137
//adding number, 5 bits max
//Varun Ved

module TestMod;
    parameter STDIN = 32'h8000_0000;

    reg [7:0] str[1:3];
    reg [4:0
