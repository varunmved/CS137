//mux4x1.v, 4x1 mulitplexor, gate synthesis
//Varun Ved

module MuxMod(s1, s0, d0, d1, d2, d3,o);
    //io
    input s0, s1, d0, d1, d2, d3;
    output o;

    //wires
    wire s0_inv,s1_inv,and0,and1,and2,and3;
    
    //build gates
    not(s0_inv,s0);
    not(s1_inv,s1);

    and(and0,d0,s0_inv,s1_inv);
    and(and1,d1,s0,s1_inv);
    and(and2,d2,s0_inv,s1);
    and(and3,d3,s0,s1);

    //or(o,and0,and1,and2,and3);
    assign o = and0 || and1 || and2 || and3;    
endmodule

module TestMod;
    
    //declare
    reg s0,s1,d0,d1,d2,d3;
    wire o;

    initial begin
        $display("Time\ts1\ts0\td0\td1\td2\td3\to");
        $display("--------------------------------");
        $monitor("%0d\t%b\t%b\t%b\t%b\t%b\t%b\t%b", $time, s1,s0, d0, d1,d2,d3, o);
    end

    initial begin
        s1= 0; s0= 0; d0= 0; d1= 0; d2= 0; d3= 0; 
		#1
		s1= 0; s0= 0; d0= 0; d1= 0; d2= 0; d3= 1; 
		#1
		s1= 0; s0= 0; d0= 0; d1= 0; d2= 1; d3= 0; 
		#1
		s1= 0; s0= 0; d0= 0; d1= 0; d2= 1; d3= 1; 
		#1
		s1= 0; s0= 0; d0= 0; d1= 1; d2= 0; d3= 0; 
		#1
		s1= 0; s0= 0; d0= 0; d1= 1; d2= 0; d3= 1; 
		#1
		s1= 0; s0= 0; d0= 0; d1= 1; d2= 1; d3= 0; 
		#1
		s1= 0; s0= 0; d0= 0; d1= 1; d2= 1; d3= 1; 
		#1
		s1= 0; s0= 0; d0= 1; d1= 0; d2= 0; d3= 0; 
		#1
		s1= 0; s0= 0; d0= 1; d1= 0; d2= 0; d3= 1; 
		#1
		s1= 0; s0= 0; d0= 1; d1= 0; d2= 1; d3= 0; 
		#1
		s1= 0; s0= 0; d0= 1; d1= 0; d2= 1; d3= 1; 
		#1
		s1= 0; s0= 0; d0= 1; d1= 1; d2= 0; d3= 0; 
		#1
		s1= 0; s0= 0; d0= 1; d1= 1; d2= 0; d3= 1; 
		#1
		s1= 0; s0= 0; d0= 1; d1= 1; d2= 1; d3= 0; 
		#1
		s1= 0; s0= 0; d0= 1; d1= 1; d2= 1; d3= 1; 
		#1
		s1= 0; s0= 1; d0= 0; d1= 0; d2= 0; d3= 0; 
		#1
		s1= 0; s0= 1; d0= 0; d1= 0; d2= 0; d3= 1; 
		#1
		s1= 0; s0= 1; d0= 0; d1= 0; d2= 1; d3= 0; 
		#1
		s1= 0; s0= 1; d0= 0; d1= 0; d2= 1; d3= 1; 
		#1
		s1= 0; s0= 1; d0= 0; d1= 1; d2= 0; d3= 0; 
		#1
		s1= 0; s0= 1; d0= 0; d1= 1; d2= 0; d3= 1; 
		#1
		s1= 0; s0= 1; d0= 0; d1= 1; d2= 1; d3= 0; 
		#1
		s1= 0; s0= 1; d0= 0; d1= 1; d2= 1; d3= 1; 
		#1
		s1= 0; s0= 1; d0= 1; d1= 0; d2= 0; d3= 0; 
		#1
		s1= 0; s0= 1; d0= 1; d1= 0; d2= 0; d3= 1; 
		#1
		s1= 0; s0= 1; d0= 1; d1= 0; d2= 1; d3= 0; 
		#1
		s1= 0; s0= 1; d0= 1; d1= 0; d2= 1; d3= 1; 
		#1
		s1= 0; s0= 1; d0= 1; d1= 1; d2= 0; d3= 0; 
		#1
		s1= 0; s0= 1; d0= 1; d1= 1; d2= 0; d3= 1; 
		#1
		s1= 0; s0= 1; d0= 1; d1= 1; d2= 1; d3= 0; 
		#1
		s1= 0; s0= 1; d0= 1; d1= 1; d2= 1; d3= 1; 
		#1
		s1= 1; s0= 0; d0= 0; d1= 0; d2= 0; d3= 0; 
		#1
		s1= 1; s0= 0; d0= 0; d1= 0; d2= 0; d3= 1; 
		#1
		s1= 1; s0= 0; d0= 0; d1= 0; d2= 1; d3= 0; 
		#1
		s1= 1; s0= 0; d0= 0; d1= 0; d2= 1; d3= 1; 
		#1
		s1= 1; s0= 0; d0= 0; d1= 1; d2= 0; d3= 0; 
		#1
		s1= 1; s0= 0; d0= 0; d1= 1; d2= 0; d3= 1; 
		#1
		s1= 1; s0= 0; d0= 0; d1= 1; d2= 1; d3= 0; 
		#1
		s1= 1; s0= 0; d0= 0; d1= 1; d2= 1; d3= 1; 
		#1
		s1= 1; s0= 0; d0= 1; d1= 0; d2= 0; d3= 0; 
		#1
		s1= 1; s0= 0; d0= 1; d1= 0; d2= 0; d3= 1; 
		#1
		s1= 1; s0= 0; d0= 1; d1= 0; d2= 1; d3= 0; 
		#1
		s1= 1; s0= 0; d0= 1; d1= 0; d2= 1; d3= 1; 
		#1
		s1= 1; s0= 0; d0= 1; d1= 1; d2= 0; d3= 0; 
		#1
		s1= 1; s0= 0; d0= 1; d1= 1; d2= 0; d3= 1; 
		#1
		s1= 1; s0= 0; d0= 1; d1= 1; d2= 1; d3= 0; 
		#1
		s1= 1; s0= 0; d0= 1; d1= 1; d2= 1; d3= 1; 
		#1
		s1= 1; s0= 1; d0= 0; d1= 0; d2= 0; d3= 0; 
		#1
		s1= 1; s0= 1; d0= 0; d1= 0; d2= 0; d3= 1; 
		#1
		s1= 1; s0= 1; d0= 0; d1= 0; d2= 1; d3= 0; 
		#1
		s1= 1; s0= 1; d0= 0; d1= 0; d2= 1; d3= 1; 
		#1
		s1= 1; s0= 1; d0= 0; d1= 1; d2= 0; d3= 0; 
		#1
		s1= 1; s0= 1; d0= 0; d1= 1; d2= 0; d3= 1; 
		#1
		s1= 1; s0= 1; d0= 0; d1= 1; d2= 1; d3= 0; 
		#1
		s1= 1; s0= 1; d0= 0; d1= 1; d2= 1; d3= 1; 
		#1
		s1= 1; s0= 1; d0= 1; d1= 0; d2= 0; d3= 0; 
		#1
		s1= 1; s0= 1; d0= 1; d1= 0; d2= 0; d3= 1; 
		#1
		s1= 1; s0= 1; d0= 1; d1= 0; d2= 1; d3= 0; 
		#1
		s1= 1; s0= 1; d0= 1; d1= 0; d2= 1; d3= 1; 
		#1
		s1= 1; s0= 1; d0= 1; d1= 1; d2= 0; d3= 0; 
		#1
		s1= 1; s0= 1; d0= 1; d1= 1; d2= 0; d3= 1; 
		#1
		s1= 1; s0= 1; d0= 1; d1= 1; d2= 1; d3= 0; 
		#1
		s1= 1; s0= 1; d0= 1; d1= 1; d2= 1; d3= 1; 
    end


endmodule
